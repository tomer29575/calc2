module
initial begin
   $display("hello calc");
   
end 
endmodule
